import top_module   :: *;

module mkTestTopMod (Empty);
	Ifc m <- topModule;
	
endmodule: mkTestTopMod
